/home/carlos/Plantillas/pruebacont/p1/cont_digito.vhd