carlos@debian.808:1587032106