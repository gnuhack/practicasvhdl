/home/carlos/Plantillas/pruebacont/p1/tb_div_frec.vhd