/home/carlos/Plantillas/pruebacont/p1/div_frec.vhd