/home/carlos/Plantillas/pruebacont/p1/tb_cont_digito.vhd